`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 30.08.2024 15:44:33
// Design Name: 
// Module Name: tb6k
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////

// Tests the pipelined_iir module for low frequency sinusoidal signal of 6kHz
// The bandstop filter should block this signal
module tb6k;

	// Inputs
	reg clk, reset;
	reg signed [31:0] x;

	// Outputs
	wire signed [31:0] y;

	// Instantiate the Unit Under Test (UUT)
	pipelined_iir uut (
		.clk(clk), 
		.reset(reset),
		.x(x), 
		.y(y)
	);

	// Generate clock with 100ns period
	initial clk = 0;
	always #50 clk = ~clk;

	// Initialize and pass sinusoidal input data of 6kHz with sampling frequency of 48kHz
	// A = [1048576, -8218189, 32107544, -81217352, 147076592, -199990256, 208937824, -168854944, 104844152, -48879952, 16314139, -3525584, 379931]
	// B = [631178, -5401947, 23050644, -63646908, 125716872, -186294288, 211911376, -186294288, 125716872, -63646908, 23050644, -5401947, 631178]
	
	initial begin
		x = 0; reset = 1; clk = 0; #100;
		reset = 1; #200;
		reset = 0; 
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
			x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;
		x = 741455; #100;
		x = 1048576; #100;
		x = 741455; #100;
		x = 0; #100;
		x = -741455; #100;
		x = -1048576; #100;
		x = -741455; #100;
		x = 0; #100;

	end
      
endmodule